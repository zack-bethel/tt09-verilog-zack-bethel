/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_lif_ZB_copy (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
  // assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  assign uio_out [6:0] = 0;
  assign uio_oe  = 1;

  // List all unused inputs to prevent warnings
  wire _unused = &{ena, clk, rst_n, 1'b0};
  // wire _unused = &{ena, uio_out, uio_oe, 1'b0};

  //instantiate LIF neuron
  lif lif1 (.current(ui_in),.clk (clk), .reset_n(rst_n) , .state(uo_out), .spike(uio_out[7]));
  // lif lif2 (.current({uio_out[7], 7'b00000000}),.clk (clk), .reset_n(rst_n) , .state(uo_out), .spike(uio_out[7])); // need new state and spike reg

  //instantiate Linear HH neuron
  // LinearHodgkinHuxleyModel HH1 (.clock(clk), .reset(rst_n), .current_in(ui_in), .dt(uio_in), .data_out(uo_out));

endmodule
